// NiosSoC_tb.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module NiosSoC_tb (
	);

	wire         niossoc_inst_mm_bridge_0_m0_waitrequest;   // NiosSoC_inst_mm_bridge_0_m0_bfm:avs_waitrequest -> NiosSoC_inst:mm_bridge_0_m0_waitrequest
	wire  [31:0] niossoc_inst_mm_bridge_0_m0_readdata;      // NiosSoC_inst_mm_bridge_0_m0_bfm:avs_readdata -> NiosSoC_inst:mm_bridge_0_m0_readdata
	wire         niossoc_inst_mm_bridge_0_m0_debugaccess;   // NiosSoC_inst:mm_bridge_0_m0_debugaccess -> NiosSoC_inst_mm_bridge_0_m0_bfm:avs_debugaccess
	wire   [9:0] niossoc_inst_mm_bridge_0_m0_address;       // NiosSoC_inst:mm_bridge_0_m0_address -> NiosSoC_inst_mm_bridge_0_m0_bfm:avs_address
	wire         niossoc_inst_mm_bridge_0_m0_read;          // NiosSoC_inst:mm_bridge_0_m0_read -> NiosSoC_inst_mm_bridge_0_m0_bfm:avs_read
	wire   [3:0] niossoc_inst_mm_bridge_0_m0_byteenable;    // NiosSoC_inst:mm_bridge_0_m0_byteenable -> NiosSoC_inst_mm_bridge_0_m0_bfm:avs_byteenable
	wire         niossoc_inst_mm_bridge_0_m0_readdatavalid; // NiosSoC_inst_mm_bridge_0_m0_bfm:avs_readdatavalid -> NiosSoC_inst:mm_bridge_0_m0_readdatavalid
	wire  [31:0] niossoc_inst_mm_bridge_0_m0_writedata;     // NiosSoC_inst:mm_bridge_0_m0_writedata -> NiosSoC_inst_mm_bridge_0_m0_bfm:avs_writedata
	wire         niossoc_inst_mm_bridge_0_m0_write;         // NiosSoC_inst:mm_bridge_0_m0_write -> NiosSoC_inst_mm_bridge_0_m0_bfm:avs_write
	wire   [0:0] niossoc_inst_mm_bridge_0_m0_burstcount;    // NiosSoC_inst:mm_bridge_0_m0_burstcount -> NiosSoC_inst_mm_bridge_0_m0_bfm:avs_burstcount
	wire         niossoc_inst_clk_bfm_clk_clk;              // NiosSoC_inst_clk_bfm:clk -> [NiosSoC_inst:clk_clk, NiosSoC_inst_mm_bridge_0_m0_bfm:clk, NiosSoC_inst_reset_bfm:clk]
	wire         niossoc_inst_reset_bfm_reset_reset;        // NiosSoC_inst_reset_bfm:reset -> [NiosSoC_inst:reset_reset_n, NiosSoC_inst_mm_bridge_0_m0_bfm:reset]

	NiosSoC niossoc_inst (
		.clk_clk                      (niossoc_inst_clk_bfm_clk_clk),              //            clk.clk
		.mm_bridge_0_m0_waitrequest   (niossoc_inst_mm_bridge_0_m0_waitrequest),   // mm_bridge_0_m0.waitrequest
		.mm_bridge_0_m0_readdata      (niossoc_inst_mm_bridge_0_m0_readdata),      //               .readdata
		.mm_bridge_0_m0_readdatavalid (niossoc_inst_mm_bridge_0_m0_readdatavalid), //               .readdatavalid
		.mm_bridge_0_m0_burstcount    (niossoc_inst_mm_bridge_0_m0_burstcount),    //               .burstcount
		.mm_bridge_0_m0_writedata     (niossoc_inst_mm_bridge_0_m0_writedata),     //               .writedata
		.mm_bridge_0_m0_address       (niossoc_inst_mm_bridge_0_m0_address),       //               .address
		.mm_bridge_0_m0_write         (niossoc_inst_mm_bridge_0_m0_write),         //               .write
		.mm_bridge_0_m0_read          (niossoc_inst_mm_bridge_0_m0_read),          //               .read
		.mm_bridge_0_m0_byteenable    (niossoc_inst_mm_bridge_0_m0_byteenable),    //               .byteenable
		.mm_bridge_0_m0_debugaccess   (niossoc_inst_mm_bridge_0_m0_debugaccess),   //               .debugaccess
		.reset_reset_n                (niossoc_inst_reset_bfm_reset_reset)         //          reset.reset_n
	);
reg vaild;
always @(posedge niossoc_inst_clk_bfm_clk_clk or negedge niossoc_inst_reset_bfm_reset_reset)
	if (!niossoc_inst_reset_bfm_reset_reset) vaild <= 1'b0;
	 else vaild <= niossoc_inst_mm_bridge_0_m0_read;
	 
assign niossoc_inst_mm_bridge_0_m0_readdatavalid = vaild;	 
assign niossoc_inst_mm_bridge_0_m0_readdata = 32'h00000000;
assign niossoc_inst_mm_bridge_0_m0_waitrequest = 1'b0;
	
	
	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) niossoc_inst_clk_bfm (
		.clk (niossoc_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_mm_slave_bfm #(
		.AV_ADDRESS_W               (10),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (1),
		.AV_WRITERESPONSE_W         (1),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (1),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (64),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) niossoc_inst_mm_bridge_0_m0_bfm (
		.clk                      (niossoc_inst_clk_bfm_clk_clk),              //       clk.clk
		.reset                    (~niossoc_inst_reset_bfm_reset_reset),       // clk_reset.reset
		.avs_writedata            (niossoc_inst_mm_bridge_0_m0_writedata),     //        s0.writedata
		.avs_burstcount           (niossoc_inst_mm_bridge_0_m0_burstcount),    //          .burstcount
		.avs_readdata             (),//niossoc_inst_mm_bridge_0_m0_readdata),      //          .readdata
		.avs_address              (niossoc_inst_mm_bridge_0_m0_address),       //          .address
		.avs_waitrequest          (),//niossoc_inst_mm_bridge_0_m0_waitrequest),   //          .waitrequest
		.avs_write                (niossoc_inst_mm_bridge_0_m0_write),         //          .write
		.avs_read                 (niossoc_inst_mm_bridge_0_m0_read),          //          .read
		.avs_byteenable           (niossoc_inst_mm_bridge_0_m0_byteenable),    //          .byteenable
		.avs_readdatavalid        (),//niossoc_inst_mm_bridge_0_m0_readdatavalid), //          .readdatavalid
		.avs_debugaccess          (niossoc_inst_mm_bridge_0_m0_debugaccess),   //          .debugaccess
		.avs_begintransfer        (1'b0),                                      // (terminated)
		.avs_beginbursttransfer   (1'b0),                                      // (terminated)
		.avs_arbiterlock          (1'b0),                                      // (terminated)
		.avs_lock                 (1'b0),                                      // (terminated)
		.avs_transactionid        (8'b00000000),                               // (terminated)
		.avs_readid               (),                                          // (terminated)
		.avs_writeid              (),                                          // (terminated)
		.avs_clken                (1'b1),                                      // (terminated)
		.avs_response             (),                                          // (terminated)
		.avs_writeresponserequest (1'b0),                                      // (terminated)
		.avs_writeresponsevalid   (),                                          // (terminated)
		.avs_readresponse         (),                                          // (terminated)
		.avs_writeresponse        ()                                           // (terminated)
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) niossoc_inst_reset_bfm (
		.reset (niossoc_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (niossoc_inst_clk_bfm_clk_clk)        //   clk.clk
	);
	
reg rstn;
initial begin 
rstn = 1'b0;
#1000;
rstn = 1'b1;
end	
wire SCLK;
wire MOSI;
wire MISO;
wire SS_n;	

wire 		     [1:0]		KEY = {1'b0,rstn};
wire 		    [33:0]		GPIO_0;
wire 		    [33:0]		GPIO_1;
//wire 		    [33:0]		GPIO_0 = {{30{1'b0}},SS_n,MISO,MOSI,SCLK};
//wire 		    [33:0]		GPIO_1 = {{30{1'b0}},SS_n,MISO,MOSI,SCLK};

assign SCLK = GPIO_0[0];	
assign MOSI = GPIO_0[1];	
assign GPIO_0[2] = MISO;	
assign SS_n = GPIO_0[3];	

assign GPIO_1[0] = SCLK;	
assign GPIO_1[1] = MOSI;
assign MISO = GPIO_1[2];
assign GPIO_1[3] = SS_n;
	

DE0_Nano DE0_Nano_inst(
	.CLOCK_50(niossoc_inst_clk_bfm_clk_clk),
	.KEY     (KEY),
	.GPIO_0  (GPIO_0),
	.GPIO_1  (GPIO_1)
);
	
endmodule
